/*
    @Copyright HIT team
    The definition of the parameters
*/
`ifndef _MACRO_VH_

`define PINS(p, len)    (p)+:(len)
`define N(n)            [(n)-1:0]
`define ZERO(n)         {(n){1'b0}}

`endif