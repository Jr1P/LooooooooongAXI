/*
    @Copyright HIT team
    The definition of the parameters in CP0
*/
`ifndef PARAMETER_TLB_VH


`define RstEnable   1
`define WriteEnable 1


`endif