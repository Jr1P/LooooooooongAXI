`timescale 1ns/100ps

// * 预解码 pre-decode
module pd (
    input [31:0] inst,

    output j
);
    
    

endmodule