`timescale 1ns/1ps

module tlb(

);

   
endmodule