/*
    @Copyright HIT team
    The definition of the Interface
*/
`ifndef INTERFACE_VH
//AXI



//Sram-Like
`define SRAM_SIZE_WIDTH 2
`define SRAM_ADDR_WIDTH 32
`define SRAM_WDATA_WIDTH 32
`define SRAM_RDATA_WIDTH 32




`endif



