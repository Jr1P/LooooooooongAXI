



`ifndef AXIHEADERS_VH
`define AXI_ID_WITH 8


`endif